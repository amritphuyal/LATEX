LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY q3 IS PORT (
	X1, X2, X3 : IN STD_LOGIC;
	F : OUT STD_LOGIC
);
END q3;

ARCHITECTURE dataflow OF q3 IS
BEGIN
	F <= (X1 AND X2 AND NOT X3) OR (X3 AND (X1 XOR X2));
END dataflow;