LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY q4_pos IS PORT (
	X1, X2, X3, X4 : IN STD_LOGIC;
	Y : OUT STD_LOGIC
);
END q4_pos;

ARCHITECTURE dataflow OF q4_pos IS

BEGIN
	Y <= (X3 OR NOT X4) AND (X2 OR X3) AND (NOT X1 OR NOT X2 OR NOT X4);
END dataflow;