LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY q5_mux2_1 IS PORT (
	S, X1, X2 : IN STD_LOGIC;
	Y : OUT STD_LOGIC
);
END q5_mux2_1;

ARCHITECTURE behavioral OF q5_mux2_1 IS
BEGIN

	PROCESS (S, X1, X2)
	BEGIN
		IF ((NOT S AND X1) OR (S AND X2)) = '1' THEN
			Y <= '1';
		ELSE
			Y <= '0';
		END IF;
	END PROCESS;
END behavioral;