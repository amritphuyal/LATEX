LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY q4_sop IS PORT (
	X1, X2, X3, X4 : IN STD_LOGIC;
	Y : OUT STD_LOGIC
);
END q4_sop;

ARCHITECTURE behavorial OF q4_sop IS
	SIGNAL Y1, Y2, Y3 : STD_LOGIC;

BEGIN

	PROCESS (X1, X2, X3, X4, Y1, Y2, Y3)

	BEGIN
		Y1 <= NOT X1 AND NOT X3;
		Y2 <= NOT X2 AND NOT X3;
		Y3 <= X1 AND X2 AND X3;
		Y <= Y1 OR Y2 OR Y3;

	END PROCESS;

END behavorial;