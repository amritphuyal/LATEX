LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY q4_sop IS PORT (
	X1, X2, X3, X4 : IN STD_LOGIC;
	Y : OUT STD_LOGIC
);
END q4_sop;

ARCHITECTURE dataflow OF q4_sop IS

BEGIN
	Y <= (NOT X1 AND NOT X3) OR (NOT X2 AND NOT X3) OR (X1 AND X2 AND X3);
END dataflow;