LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY q4_pos IS PORT (
	X1, X2, X3, X4 : IN STD_LOGIC;
	Y : OUT STD_LOGIC
);
END q4_pos;

ARCHITECTURE behavorial OF q4_pos IS
	SIGNAL Y1, Y2, Y3 : STD_LOGIC;

BEGIN

	PROCESS (X1, X2, X3, X4, Y1, Y2, Y3)

	BEGIN
		Y1 <= X3 OR NOT X4;
		Y2 <= X2 OR X3;
		Y3 <= NOT X1 OR NOT X2 OR NOT X4;
		Y <= Y1 AND Y2 AND Y3;

	END PROCESS;

END behavorial;